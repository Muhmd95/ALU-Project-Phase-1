module ALU_Top (
    input  [9:0] SW,   // The 10 Switches on the board
    output [9:0] LEDR  // The 10 Red LEDs on the board
);

    // TODO: Declare wires to split SW into A, B, and OpCode

    // TODO: Instantiate your ALU_Core here

    // TODO: Connect the ALU output to LEDR

endmodule