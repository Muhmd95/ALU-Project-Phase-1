`timescale 1ns / 1ps

module ALU_tb;

    // TODO: Declare registers for Inputs (reg)
    // TODO: Declare wires for Outputs (wire)

    // TODO: Instantiate the Unit Under Test (ALU_Core)

    initial begin
        // TODO: Write your test cases here
        // e.g., A = 2; B = 3; OpCode = 0; #10;
    end

endmodule